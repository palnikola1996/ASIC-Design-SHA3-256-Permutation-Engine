parameter X = 5;
parameter Y = 5;
parameter Z = 64;

parameter RC_00   = 64'h0000000000000001;	parameter RC_03   = 64'h8000000080008000;	parameter RC_06   = 64'h8000000080008081;	parameter RC_09   = 64'h0000000000000088;	
parameter RC_01   = 64'h0000000000008082;	parameter RC_04   = 64'h000000000000808B;	parameter RC_07   = 64'h8000000000008009;	parameter RC_10   = 64'h0000000080008009;	
parameter RC_02   = 64'h800000000000808A;	parameter RC_05   = 64'h0000000080000001;	parameter RC_08   = 64'h000000000000008A;	parameter RC_11   = 64'h000000008000000A;

parameter RC_12   = 64'h000000008000808B;   parameter RC_15   = 64'h8000000000008003;   parameter RC_18   = 64'h000000000000800A;   parameter RC_21   = 64'h8000000000008080;
parameter RC_13   = 64'h800000000000008B;   parameter RC_16   = 64'h8000000000008002;   parameter RC_19   = 64'h800000008000000A;   parameter RC_22   = 64'h0000000080000001;
parameter RC_14   = 64'h8000000000008089;   parameter RC_17   = 64'h8000000000000080;   parameter RC_20   = 64'h8000000080008081;   parameter RC_23   = 64'h8000000080008008;
