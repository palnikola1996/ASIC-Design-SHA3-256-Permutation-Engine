`include "./theta.sv"
`include "./rho.sv"
`include "./pie.sv"
`include "./chi.sv"
`include "./iota.sv"
`include "./permutation.sv"
`include "./string2array.sv"
`include "./array2string.sv"
`include "./pipeline.sv"
